module ro_gen_0 (
  input  wire en,
  output wire y
);


INV_X2P5M_A9TH  u_inv_DONT_TOUCH_inst0 (.A (y_inv_dly), .Y(y_inv0));
INV_X2P5M_A9TH  u_inv_DONT_TOUCH_inst1 (.A (y_inv0),    .Y(y_inv1));
INV_X2P5M_A9TH  u_inv_DONT_TOUCH_inst2 (.A (y_inv1),    .Y(y_inv2));
DLY4_X0P5M_A9TH u_inv_DONT_TOUCH_dly0  (.A (y_inv2),    .Y(y_inv_dly));
assign y = en & y_inv_dly;
//A2ISO_X2M_A9TH u_iso_DONT_TOUCH_inst ( .A (y_inv_dly), .EN (en), .Y (y));

endmodule

module ro_gen_1 (
  input  wire en,
  output wire y
);


INV_X2P5M_A9TH  u_inv_DONT_TOUCH_inst0 (.A (y_inv_dly), .Y(y_inv0));
INV_X2P5M_A9TH  u_inv_DONT_TOUCH_inst1 (.A (y_inv0),    .Y(y_inv1));
INV_X2P5M_A9TH  u_inv_DONT_TOUCH_inst2 (.A (y_inv1),    .Y(y_inv2));
DLY4_X0P5M_A9TH u_inv_DONT_TOUCH_dly0  (.A (y_inv2),    .Y(y_inv_dly));
assign y = en & y_inv_dly;
//A2ISO_X2M_A9TH u_iso_DONT_TOUCH_inst ( .A (y_inv_dly), .EN (en), .Y (y));

endmodule

module ro_gen_2 (
  input  wire en,
  output wire y
);


INV_X2P5M_A9TH  u_inv_DONT_TOUCH_inst0 (.A (y_inv_dly), .Y(y_inv0));
INV_X2P5M_A9TH  u_inv_DONT_TOUCH_inst1 (.A (y_inv0),    .Y(y_inv1));
INV_X2P5M_A9TH  u_inv_DONT_TOUCH_inst2 (.A (y_inv1),    .Y(y_inv2));
DLY4_X0P5M_A9TH u_inv_DONT_TOUCH_dly0  (.A (y_inv2),    .Y(y_inv_dly));
assign y = en & y_inv_dly;
//A2ISO_X2M_A9TH u_iso_DONT_TOUCH_inst ( .A (y_inv_dly), .EN (en), .Y (y));

endmodule

module ro_gen_3 (
  input  wire en,
  output wire y
);


INV_X2P5M_A9TH  u_inv_DONT_TOUCH_inst0 (.A (y_inv_dly), .Y(y_inv0));
INV_X2P5M_A9TH  u_inv_DONT_TOUCH_inst1 (.A (y_inv0),    .Y(y_inv1));
INV_X2P5M_A9TH  u_inv_DONT_TOUCH_inst2 (.A (y_inv1),    .Y(y_inv2));
DLY4_X0P5M_A9TH u_inv_DONT_TOUCH_dly0  (.A (y_inv2),    .Y(y_inv_dly));
assign y = en & y_inv_dly;
//A2ISO_X2M_A9TH u_iso_DONT_TOUCH_inst ( .A (y_inv_dly), .EN (en), .Y (y));

endmodule

module ro_gen_4 (
  input  wire en,
  output wire y
);


INV_X2P5M_A9TH  u_inv_DONT_TOUCH_inst0 (.A (y_inv_dly), .Y(y_inv0));
INV_X2P5M_A9TH  u_inv_DONT_TOUCH_inst1 (.A (y_inv0),    .Y(y_inv1));
INV_X2P5M_A9TH  u_inv_DONT_TOUCH_inst2 (.A (y_inv1),    .Y(y_inv2));
DLY4_X0P5M_A9TH u_inv_DONT_TOUCH_dly0  (.A (y_inv2),    .Y(y_inv_dly));
assign y = en & y_inv_dly;
//A2ISO_X2M_A9TH u_iso_DONT_TOUCH_inst ( .A (y_inv_dly), .EN (en), .Y (y));

endmodule

module ro_gen_5 (
  input  wire en,
  output wire y
);


INV_X2P5M_A9TH  u_inv_DONT_TOUCH_inst0 (.A (y_inv_dly), .Y(y_inv0));
INV_X2P5M_A9TH  u_inv_DONT_TOUCH_inst1 (.A (y_inv0),    .Y(y_inv1));
INV_X2P5M_A9TH  u_inv_DONT_TOUCH_inst2 (.A (y_inv1),    .Y(y_inv2));
DLY4_X0P5M_A9TH u_inv_DONT_TOUCH_dly0  (.A (y_inv2),    .Y(y_inv_dly));
assign y = en & y_inv_dly;
//A2ISO_X2M_A9TH u_iso_DONT_TOUCH_inst ( .A (y_inv_dly), .EN (en), .Y (y));

endmodule

module ro_gen_6 (
  input  wire en,
  output wire y
);


INV_X2P5M_A9TH  u_inv_DONT_TOUCH_inst0 (.A (y_inv_dly), .Y(y_inv0));
INV_X2P5M_A9TH  u_inv_DONT_TOUCH_inst1 (.A (y_inv0),    .Y(y_inv1));
INV_X2P5M_A9TH  u_inv_DONT_TOUCH_inst2 (.A (y_inv1),    .Y(y_inv2));
DLY4_X0P5M_A9TH u_inv_DONT_TOUCH_dly0  (.A (y_inv2),    .Y(y_inv_dly));
assign y = en & y_inv_dly;
//A2ISO_X2M_A9TH u_iso_DONT_TOUCH_inst ( .A (y_inv_dly), .EN (en), .Y (y));

endmodule

module ro_gen_7 (
  input  wire en,
  output wire y
);


INV_X2P5M_A9TH  u_inv_DONT_TOUCH_inst0 (.A (y_inv_dly), .Y(y_inv0));
INV_X2P5M_A9TH  u_inv_DONT_TOUCH_inst1 (.A (y_inv0),    .Y(y_inv1));
INV_X2P5M_A9TH  u_inv_DONT_TOUCH_inst2 (.A (y_inv1),    .Y(y_inv2));
DLY4_X0P5M_A9TH u_inv_DONT_TOUCH_dly0  (.A (y_inv2),    .Y(y_inv_dly));
assign y = en & y_inv_dly;
//A2ISO_X2M_A9TH u_iso_DONT_TOUCH_inst ( .A (y_inv_dly), .EN (en), .Y (y));

endmodule

